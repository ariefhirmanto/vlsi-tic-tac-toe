module controlunit();
    