module q_accelerator();
